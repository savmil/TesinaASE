--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:12:59 11/12/2017
-- Design Name:   
-- Module Name:   /home/sav/ASE/gestore_display/gestore_display_testbench.vhd
-- Project Name:  gestore_display
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: gestore_display
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY gestore_display_testbench IS
END gestore_display_testbench;
 
ARCHITECTURE behavior OF gestore_display_testbench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT gestore_display
    PORT(
			number: in STD_LOGIC_VECTOR(15 downto 0);
         enable : IN  std_logic;
         clk : IN  std_logic;
			point: IN std_logic_vector(3 downto 0);
         reset : IN  std_logic;
         anode : OUT  std_logic_vector(3 downto 0);
         cathode : OUT  std_logic_vector(6 downto 0)
        );
    END COMPONENT;
    

   --Inputs
	signal number : std_logic_vector(15 downto 0):=(others=>'0');
   signal enable : std_logic := '0';
   signal clk : std_logic := '0';
	signal point : std_logic_vector (3 downto 0 ) :=(others=>'0');
   signal reset : std_logic := '0';
 	--Outputs
   signal anode : std_logic_vector(3 downto 0);
   signal cathode : std_logic_vector(6 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: gestore_display PORT MAP (
			 number=>number,
          enable => enable,
          clk => clk,
			 point=>point,
          reset => reset,
          anode => anode,
          cathode => cathode
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		reset<='1';
		enable<='1';
		number<="0000111100001111";
		wait for 10 ns;

      -- insert stimulus here 

      wait;
   end process;

END;
