XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~�A"�����'�� ���/�:�D���T��N�
f0�h9�]�o�+x�w���h���O4;�p���Z��l�L�g/L�fv`������bL�`�t�Bm�2�M*�����)=5&������~�QS���y��@�?d�N��$�ys7.��� ��{����r� ���9'K�5qJT��=���ҽ7��)H�%�V8hJH��:E?o�c46���k���3�2���Bő���,u��M�4��Kټi��"��װ��p����_ &�G���^}x ��z�
O�[h��Ah3����X|������l� �笢��SW��[_o#���=����6I�e�(Й�`\�{��{�@�7/c�4 ��ǀ���S��ǄcîJ����XfM�-
o�
q4|/X�.�V��\i��N�	Z���	(cZO�j=�rX��<jE�iU
�|غo���٦��,na�2[p�w�攙~+O�~��B�"W�!�ĸs�M����W�f Gs� �9v���]3!ݸ-?-5�Q��0��Z�D��B,�C_�vg3�o�_>�d0\k$�jh�kD�P�c�b3 ���_�¯����E��@���#fQ=��h��7%���� �Я�Ċ]���Y���!{����0�ڐ[%�*�g�F�;��AV��a�����>��j9�=�sw��_<���Ƭ��3�|�ױM�X�k-�^x�J�r1�\E�򏷨Ш�b����qx��RTC�B�*�XlxVHYEB    3189     890�f���������v�1ůc:M}�M��[͕�?Gk-瑜e� �q3yhlT�&�h��GW��.�t����q�-5*L"&��(ۻ�$C�����,/+��X(4��wE>9��݂ͩߕʁk�ZW��"e�J��w��(V��GBR���T~ h���L�`0??(��rM�/7�s}�6.C��A�\���굱�k�<����oD�j�[T�� U_4i������.��KMS��,���7����>��l��1rml�h�S��Z���B�[�Zf:��Xw�۴����>�4�d0փ?�-+XW��7�\����&{�������,��TFje�Wb�}�p�ܣ�����^�acf@vG�fm�XA�8��a��6� =����`�^I.@�0�1��V~HP:$0p�ޓ�) %��)șo»=L���O���7'W�AG2�#�V�d/��1�ن�W�,P�x}�o�w��3b:־���XR< h5k:�(�W����k��*��I ��I��&:�h�s���bE�є���?$�Jx �l'�lo��;훯%#;v�ˈ�
~�犈;��vvd����O�T��o��L�T�y��]�P�>)���O�ǐs?}�%�#w��e��+��o�$���D��P7����)���t��!�b2F���fw�~��y3o�ʮ<R���5⋚8j
���sK�8��"�,��ͯQz�i�[08�W�@��<�Տ[7?]E�z�٥Q!�1L5g�l&��a��HX�b�\��h)d�2�K*З� �IE�J/��<�v>;�6@J��g2tw���ME��@���#Cm9Q_ .6S���.�B��s��;A�s�`o�I�x��� 4&���-w����"�Bн����R~]���(V 9K��]���b��"O����[�Z��&5��#���a:�E��a�M4` ځeO�Wp�ڍ��YQKy�;��({M.�G�S�G�s�3���T�{w#�����!�k�ԛ	���-x��TA-w�"�����g��j�s�&}���;�������V(2�����̬1�#��+�u#�b�cqd��/�����jK�h6tU���7~]?n��ren4�@֬"��g������P�Ru�3�r���f��sEf��ؚVlx>m�o2���T���Յ>q")e�b2o����i����-Q��7|�ȱ%��o뷝L.��D�K�o7Ϛ{3�����|󩵡S���0��k���%�u�|Z6��qj��k��V�qF=�V���{�7������&a:���s��3K�AcA��iq�<��b�}�t%6�l�U7u? ����7������+�`Ň��g+���s���A�Wt3 h$6�(m�5���C�9q�c��{u�r��>Zȧ��ZR��p@�i�pQ�ٟp�fo�&I���H�D��(j�0bq-Z����LŘ��7�E~���Kj�y�g�ہ6"u�r�7�� %d��m�5�ll~��{�]����+��G��g98JT7�f�7J�9�ċ�q��zI���4�\��=�T9�5�۔�
C�y���s���.�aixb��x���1/��H��A`pµ)0��~�W俌��Xm�,*2�+RZ0�&ɴ@��5��8�3�r�aa&�&ߏ��a�����~ 
��~�i��{��tI�ݙ_�A�(̂�p�uN%���W�iy�V�GQ;��!�E("�
B	c|b��h{
%�2���G.��R.�f_�Iۃ�k\bi�E]wԮ���x��4�И�BB�k�U�ا�l2��� ��E�Xg{�TN��$�nΩ��G�լM`�̗cl�qcR���q����> Ч����vyx/���HYp�.*�\Y��P-�2$���� �8�n��O�;j���a�%�-��M$	�D�f�J��肤�R�	�Iɻ^�F$ed�m�׳���.��q�r�ڴ
_'K����[¤n�/��X`�Ӛ�.ݗ��\k_.W\>f?�oiq�V�-�D2`�{�X��kvb}p�[��ǖ'��E�4��A~B.~��&	�Wġ�#y_���c���>$�H;��)�'��Z�ljy�����6�*�-G*�-}s�m���N\�<^�;H�g!�t�7���C� e=�Ռ