XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o�/Z��8��
:uo�)K���(}?h�6JӦlo0���0�p�����زj�w0��7`���X�DA/��!i�g�}�u�y��Y�.{���W�n�vLZG]�����$Ӗk�!�f��/RT���W ��<�$x�L�Fk}�X�[l�-�Х�1�^�y%��s�C���*y'�؛�H�<���Js��+lB�M��u��p&�I�>ƻx����띈�oh�s_%3��Z,&�S��YFͻ�`���p��wD69���	��f?5
��$@��$$�;\4*���P�G�J�I���h�v���6����W]��Q���}�U���f2M&��(��n������Cj����=^͢,<A����>m�>�
�p0�P�!8^g}o��㵀��tWpu���d�B�"��bU�;�$��#z�h�-u��Iɢ�����m�����s\I�=Py:o�	jOM��Mm<��.Ch����9x�"�)Uf��� ~"2|Di��Cc0�8g/i���̒e}<j�w�`|gh��,g����W���������Ş��M���Y�{n^����P�Zf|F<�:ݍ^r܂�0���U��f��� T3.����W���~�]�ؙ��"��εj��������EB\�a�'&��7��c񨓠�U�V�������ە>W��z	Պ�����3��RDp\���BF� 6��eXY��׾�����X�R�."��D�eù2����jH�:�ˣ@����@��A��һXlxVHYEB    5ee8    14d0���
ƺ_"$��f�[��`�ҝ��b�G������4۞p%�盛W�̨��0��#`�4�n���]y���	���T2��I���}.c��nak.�j9��_1?ob|��m�gJ�9��g^�ݞ�T}�0H��xDs ���(�I5pZ>(���E��I��ϻ.9����y5/�1��# ����r��n�"�@v^��z0Y�k=ϞmB*UO�K.|ޜ�~�S�z-Ncj��=v�}��=M诐L�ʛA�z&W�Q�x~a� �g��M�`@q��y��H���� C��	��R�Y�_ s�$�n$I�Ŵ0�b����9�:����{�TM���.����S[�O���ص�����}�L���T�X�{8"����FI�$�F��K^�W�[ȏ𐐮��p(Tv�?�m��3FBp����\s^A�.�T�O�V��@��j-��^@��&�j�����/�g��E]�����-ëq	8����/� ��#�*C�Ph�`�Sh��Е�zݘ//l��9�8u#w$�vb�L��~�Q����,/L�.�FcE��x-�lbWeqMO��)ó*��$v%�vMȸ,T^M\�)�&�l��b�qW�~�Ka����P�$GeP~[�e�4,������}�"V�Etn�ʫ��q�[�&��o��$�ؾ@�>:��t���q�>:��9��B7���d�m�]K��\2]@�$�M]\
�~,p�C��6��a�j��̳��>�uac7�1�邤i��l���D U0%z$�/o���.�q��F�0�M�Η/|���A_�C�Z��;�6{ȾZ���3N�v�x<�s1���<U�67�tl]��=���CΫv^l�_���!��Ρ׳�� 	��q�H�F�/5���^����h��� �iQ�rP��7�٧e��+z/�oa�����&���������g��W�^�
YL&��B}4�Te�ly1�b�n�Ln
yy�% g]��P]�n�����>��.fP�tZ�<�Yq.�W��í�p�B_�E܄��һ���T�r@��,��Q��)�]�"�xjb#�o�Ń��I������!w�l�E���$�(6d�@Z�[d���)�����	���a4';���
+ݞ�-���H�s�dͤI�� 5́#S0�O��{�PQӢ_	3���a��4S�~Ȥ���q����I&6�G�$HZ�p3��25.��Ew+�,�?kQ�)i=�?n`�J��$wM,x/@����퍘�qu��ou�"��+Uc��9�Ev=�Q���M.AW�L�+�5�8�4Pp�O����b����e���k ��ߢ����U��]-��޴D�*�;���*��gQ{miD���l<ނ��JS[�KqL!�zX$�����w"�4w��o��9B$҂I/8pm	�5��KY�6���
>ئ�
+b���w�,9��f�F�ƶ��ȁZpT��Kvy� �9G���a�5b�H��,Q"�X�Į�g����|U4K�.s��%�s�+��__v�r��Ɓ��l'�si*H���E��	�<�ha�ًN�d�� ЅgK��+δ��l�~�����q�<���IE����>���k��<��,��C�g[x����;xĴrz�Hj]G��*�Hm�h�B7�R|\SC����Wh�=�B�~S��j��H4]R�8E)��*r�J�̧�������̩�F%e���즑oiBl�>�%3�7�"�	G�+��:a�KGx۷l�d�,p�ʕ)6$��=��"Ul����k&\�e�[&�� r*����/6z$}�I�V��^<����&�*n�ջ�
��Y)�	� �����*��v<�Ƒ��uA�DI2��=�����?d�������_���1o<��z�^�5a� ,{H<�K}��U�@�������KO?W�V�)���w�K̒m���t�[�Y�F;$���S����an��D��eCpiDcx�,�͏~g�WA1��0TB��ZzSk�K�V��֧����EĆVt7��c����������i��thGJ��+Xpkr�5t	��<հK��������fLY},?Pl5L�_,��}���2���3�^�1�� vtF+�6OZ����	m0��z��Q*�z��4g��L;�@����� `r�Y���ʝ��4�"��cCͽ�l��WE�|�ɾ�`�Bj��S�j�1��BGvi��9(���!�('G���f�f4s���"S�v9*�3�!�7�Hs#�����7�Q�����R*}���b� ~�Ԝ��B���a{V��m%&[�)��ӻ��S���6#bv~�ȷS��@��,uw"[�xf�)��%��<�y�^�IAL묓�n��؇\(	RoO8�m-D��0������P�˅�%��M%�(!�)���
��(f�T�.[i��\��!T�P�0u�mR��n��U�R��8�@���5�8�I��>q{�V9���G��Mz����bn�z�z��ЅI=Ν� e�f��G�i���^V�ǐ�q���!5o8�m�<�6e<"O`�D��3�ˀ+[��&�w��D�ߗo�tr�ti}��D�N��O[��)k�Yȗ	��Db�~�-�]#IC`�u�|D���֥�wv�\ -9�T��L��|C�V��ߞ�3�U8����;�?f 8�|��B�-"!����,F��k��r�����9�6M�ސ�pr����ʌ�B&"��wV$���!Ĉ�1v#a4�����ɕ٥�=�^w�:�޲�Y~�u��%�A��C{�9Qh��'C����	�k7��~�CMh�W��ƎU��=O7p�SV��޷ј����<4���f��}�4d�Z�α�V�Pлڱɦ�w�&������D�	SJ`G�@�e_䩏�'p���AX���Ɔ���;��G8�ާ�dŲ:b`rk��oϺV3o��g~��IΑ�G�	 �<�����׫�7�_!w:�(q̈́E�IW�I�?Ƭ���D�{�*Y�<.�]s77��e���Miְh/g�R�-l_�̷��9ηZ��#�_�[��Q��b0�3�s�G,�(����2�e�߳_e���~��Φ�X��ל,��Ih#�H3��vA�a�ѹ_Έ��S��z��L���1`�*L�ҕ�6a�#i9�;��9p�l�O�;�T�W���(Y��>Λ�!�'��"~H*�^t8� ��
q��gz{�,�		�b	&+��^/Z�J=Qy����>�e���xc�|�Ms���!����_��>�MCX=�C��ՕT�4���ۿ�Sy�WUx������Y	�fU�z�fNU�~���DZ���#�6��,�b��ui$�(�=�>�dHo?�����ڊb�����Β$Է����l�j4�gf�xz�(l������ˉ�>rZ����X)`��Ҍ�y[�D�+U6��	�=��q�WY_2�?�4w�1&�W����$D���bL��\T��Ә��|�ʹyj�k�TQ��G��g����$����U��h�ʤ�K��]r�v��Y��t�Qc^=U�4���9zB6��^UA>���.�i}�S���c���b�h-i-H��G��'�5��9��O�ӡ�`��<e8߬��t��vTHu �2��@K�1`�3ٕ�f��w��mt���r���KM+�cA�ns�J��@^�z�f͖"gP
��Lq�����E�%��kz5�q�=�B6W�(hJ�
f�O�y�%�<���=��>��l�RZc]��H�=jz����d(�]*�&dr.>rxy�u*i,R���i%h�P؄��}/}w�<j`a����>�*�5��b�7�B���t}�����M���
��h��~�=���p�}@���n"$��Rz�E��7��-�v���0tI���x+���T�ߧ����s�E�F��y��/mڀ�d�a�d?O쓰)*U뱚��;�VH6�t��'�x���ht;3�~�%��%�A�pl��_e�\��)��)��(dJ:�D�!{�1�� 5=mզ+���s#�_$dx	��@�QC}-�@uc������Xfi�aJ?AI�R��,��p�2�ȸ"]�Q�g�)N���9~���`��D��2x��{zC�'�=k����Jlu�j"��Si�t��>�y��4m�ࣗqƂX:�	[9�c(LY�δ�[��/�]��,�KS����c)��j:de-um�	m_���g']������h4�v�F0�eV�?+����m�Oqv���d����� w�ɵ�ᾐ
�r��T�����i9� �j-��l���Y�C�ߗ�nLX��$E��`�沓X�� �21�$S�f��{��58���Ht�f�O���9f�u��9�w�����["9$B�D����ːa�?�A��^�izS��\X2��	�!1�Il��i�q�QʞO�{�K�l>7�:Ȼ��Yy	�4���R�Ӿ�Y������O#��U�燖;�|6�-X�vѽ.�y���:��@�������n~�Y��o�J���eZ� �G�5�(\�����4%�$��|}p��_�ef��P-�i�]��������Ҭk�sI���"J���"�
�l+����԰�z'K�K��\R#o�mX%Yt�Gc�21�(]w���ɒ>�ʕs}���_%`'TU"JL�k��MEZO�k�~�w"#-�+�{`?z�=}��Gż�Jv���Y�Н�'���<���.	� �C�Up�[�t�>�VG5S]2H�ŵV�߿�y:sU!�,��dW��g�+i����J��Iw��0RDD�?��?�z��1�5eԇ�U���y�R�s�w��>EQ��5
���Q��W���+}�u���r�B�3E�p�n�WJp���xO�H$��!@�k��6�V�z�e7d��/�)`,8<��h�Pz���Rآ%����EOv#C���q�!�2 ���;rMBU��"�nBM:����JIDHLl�ZZ=�C�����M!�fxP�G��PF���Br>_]�P2���>��E�d��C���� y����~�b}*��>a0|4ߟg�J�{k=b����64`K�~5Ý΄
�B532�a��g�K�n`���D�­��f�҇8�����C,9���h+�G4���]*�|�����6o�;�$I�=,+)�_�����M�-�
���k!̊
*�Q�g��Ei������d�