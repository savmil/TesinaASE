--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   12:35:30 11/01/2017
-- Design Name:   
-- Module Name:   C:/Users/Public/ISE/cathode_manager/cathode_encoder_testbench.vhd
-- Project Name:  cathode_manager
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cathode_encoder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

ENTITY cathode_encoder_testbench IS
END cathode_encoder_testbench;

ARCHITECTURE behavior OF cathode_encoder_testbench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cathode_encoder
    PORT(
         nibble : IN  std_logic_vector(3 downto 0);
         cathodes : OUT  std_logic_vector(6 downto 0)
--			anode : OUT std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal nibble : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal cathodes : std_logic_vector(6 downto 0);
--	signal anode : std_logic;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cathode_encoder PORT MAP (
          nibble => nibble,
          cathodes => cathodes
--			 anode => anode
        );

   -- Clock process definitions
   --<clock>_process :process
   --begin
		--<clock> <= '0';
		--wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      --wait for <clock>_period*10;

      -- insert stimulus here 
		for i in 0 to 15 loop
			nibble <= conv_std_logic_vector(i, 4);
			wait for 50 ns;
		end loop;
      wait;
   end process;

END;
