XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&��j����o'���n�L��wxP�x��@/�����	�i��CP� �5<�G�F>^ش�"�W��ڜ�A��8s�O·"E������.q�y��ێ�!GVRۄ~�Xc���\�����z[�	u�/�>^8Z'�ҕf_��ppF�t�I�8���������׮���|)��Cع�+D�5�s����IP)=��)'��]k>�E�n��5�Z�� �5G?��\  [kM���X+�`z�=�����d4.���S�����fq�!����2[�HI6�n������=x�s�+�f�p�uqKO[.X��g�;p��Xܢ�z�)�����%��\%M>,bn��F?�TB�B�.��hK��n����A%��7X�����n��˜mj��w�,@�����g�ޖ�G~��a�`^�b�\�vq"0Q����0�E�X��2���=�O&�����`f�=���ܱc:����XX�Mh�b.�i3;UGĳ<.;�p���0��B�3:ވ���M��"(��<,ԝô(0�͎\�I���A}\e�\��u0�=�o��-�ێ��B�&���&�4�RLA�a7 ��mͼ�3Js�W���҄���=fO,v��b�U����(4t�Ӟ"��hă�LwbǱ;�~�o[�͇"k����Z��Γ�d��]Hhb����?'knC���f��� �P;�O�+Dw��z� �3A�����u��7�&�@�½����C*�by�3��qYϧXlxVHYEB    1795     7b0'�DW���p�0��PD��0_n��bp��A(E�P�|�B���3sXl����w#��|��և��v'�ΣZ���H8����~Y��o�V���0�H�P����-�7IH�)��[�t4����w5�'��A��� ÿt��G#����6B�`�L� �r�C�&BБ�1J��J�C:�Q��_,�'�볤����a̯�V5�z���3[v7�����K�`ʕ�뱡cyR�5�l%��MLK�yƤ�m-Q��	Zǃ�xYOc~pj�8�����A��uz@-�e_%F@|`��W�ٓ-L�?-ǯ��p�ăE"X�v d`��~��������-d'x�S`��e��\mT�&��<I˷���st���Y��R:����:�����67$,k� ���8�t ��uNs�.�zUr���l���K_���Z�۾���Q���Y{r 쟲��V�"���Ȍ�w"��GPMLp[ �ȋC�6�p��!~V��r��r��'n�.��aT��s�J������K�����1ľ�|�XI�Qf��,�Y�4�gޑ�9�Na��Ϊ��M�*�z���9n:��W�"��>Ӵ��0u�ja���h���귲��G�ǏE>3��d��$Jw�i�6m5��?�Ꮆ�l��WL_�El�I�s�9�f�N.��H�B�O{-�1���3W22�^�%���ǧb�vA�$VY1>D�E�.�>�,d�˘����me��]���G_
���y\e���0 �j5�@	�7���`nTq�@���0*{���q��h��x3��<=�p�J���-Yܽ���Q���ٓ(�gh?i�����޵P]��8�"E��Tص�����X,��Զ�{	�
]�a�ǯ�쟠�:��!.)�} �^���ٿ|��vz��'ʤ�������{)X�o�1�i���Ov���.��t��V����"ٲll��1�>ٯ��w?b��+B|}�B{��O��뗿��;���d��Ŵ�a1���O�ڕ�<�RG�����WSZ��R��`�	��p��(7�h�w���}�6m\�[{�����̕���p���6iS��=u�� ����v�p��ޑ���[�t(3v�5q��^9̂��(�e�$���Rr�ʚ]���e���/�uW��,�ڮs�c��ys���$�����{����Z�z���,*C�4<- ��r,u���I@J���&2�d�78B����s��a��r��U��@Z2�4�� 1x8��5�m>�����nt�U9r�0�VE|��*�e�J%��" ��y��(�IX1��{&��p�&�MP�{"�S^ο>*��\%5.���O �@z�凜�*S�S)�P-����ak�yk8�k��kR[=d���oQݭF���R�IU�O�W�(��ѭM��� �?Knΐ�F� qL�G���u���dɏ�ZÅ��Pl�ds����!K�O�U'����?�����}(�8�U_��r�ԛ�tܩ;��z�<^.��m�x�`�[��&�����ۘvtB�@��&��qȗӧ���g҅�KY�Ah>�g��(	ܖw%^����;��9L�Bk��&��2��I��<��lR���[�kW
�NǏ�hf[R���!yQ�(��^I��J^uR�G���(>�t��\������6l���-��L���F�UX�tM���`�us���z�1Ɔ�)��V�!ʙD��`�a+ɶ_�B|�V{��I�t�h�P��<�}���o�A8�W�s�
Q�9%�P%Z����b�Ԩ�\2G�}^����*�&x����<����+�v�>W�U���|�nP�a휊�{}�0Ɯ{0ÁF���IqL]�D����R����l>Z�'��e(��?l��n���8u������QK�@p�bP݉�iOl6���B���_��:�