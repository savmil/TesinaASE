XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����/m�`�@ 2n�K���:{:_�_��	G
�#DL�¤���?�d9�*RP�|��x��v;�)4��V*N���=��'g��Z�-TQ%f���KQ��l��T�^�kv�v��@8�7UN����)8�g}���0)/��ـ�!�t�- �\���Mu����u�A������$�u曍/ �~L�l!�;�L7� ��A@Q�m[��S�J�Sz���!(�o��드��� �-��O�V~Q����ֻ�oZsy��$2U0��&�5������rQ4��Sc�s�+�\��JVg1M��������SV�Q���(2w�o���g��Ԕ�/���������+�Y�}i2Z��|��713g�ƚ�r;�b:���گ*���$LQ
ل4��v!��& ���dj
+��7+ԃ�u�`����&?qr;O�n��d}I�����Ѥ�;!� �����M�aH��͑O�c��5��;?����0�,�<s6WZ�<y�	"��o���Z�����{Q��kD�Ȣe�]3�,{�)m�$N��Lv�y�A��5ez0j�Q�bmB�ܗ�t�����y��>/�G�"b�������'HDy��|���F1Kd b
�x�|�Pc��y�/�vC�t���2��e?J��;���S��O)`��%?ji0=)|�3����b��W
�1_����4�"*������~�f�Rv4&���yJy����<P�7-8�6^��/t�?�Sm��줲� ĭ��z��Z��I��XlxVHYEB    3357     c80H@�	h%�ٿ��T���'��%��Ũ��5����>�?;�P�4D���������d����#Ȩ��]��M������y���l@#�ఄ8`9c���/_:(���'��Sѿ��=�`����uu �`��� �sM&?�f�ӭsKnR��p�o����A����e\�������V�J��+q�(������X�D1�:�-{�yxoaUx��Ѓ|�!���d��
�	�ŭ=K�n���@6ȋ�Rȵ&�o��.���v�*cgQ7��eN�*x��y�x�%��"�a�<6hY�aQ>YV���-��0���Q�}�����yM1�̈؈�3�w�K![�GH��
�vaR7�&V�9�ʴ�?�<߸m�N2�6�͈Cp^����.!G�>F7�Q���e���d5Nk���a�ԅP��EN��o����s4c����k7��D��>ҔN���E6��L�Ɯi���=�����&�Un��\�Z�t1��šB���>�]k�C\�Vޔ�\�����K���������(���[�N��#�8��Q0���SE*���	͛�:���g,�#$��H��|�|�8h���aD�x[[W��y^�Y����^H���P<z��ƲL����,N=Q��	xi�E���%��aa[N��}�2`�tP�l�X#6�l��������B�T� ��#jfb;�ե���|�k�)t�)�V�j�I����i��5�\����ԤPE�g�+�jZ@�7����D�	v8-�$������r"��q���]-���$��Q� �(��L�wH�qDB^
�s���f��|�ŏg�E@�!����Zn�~��0�����{L��V¢���Ǿ=p�]dq�?��wϘW�;l����g��n�\�d�.�l����]�FB3�Gĕ�;��Zd[ >
8��Q,(֟F��됛�'�[���p���'l�Wuݴ�Y[���g���-zy8~}~�Br#(5�z�����>c���"y5��-��4�D�'������^}������8�o�E�L> t��5�Fh���Q�p�G��R?+AC:�����rEY2����<����繌����X'lK��{�yh|M���M�
�]G|-*�M�MXϹ���Ɖ��G~����y|p�(��˧m4�g��ut6�������)l1@艶���}�ܡ�ק0T�c��l}p?����Y������K�q�ǃg���CtJ�Fzh�	5o�޷$���<���� ɠb:�	� )�����'�mi8�>&�����T��t-�]�Q#��I�)Ɣ�M��crVIjt'�q-Ha n�@��ԛ���#=K;W�+ѷͧK�Eq^��P���vk���q��Y�	�_�oIY{.���ʹ�^�&�������r�#3�{;�XH�B��@d��[�'�~�*��p���ж�]�+�=z7�n�QS����s�l�����=e�����̧���3�qV�~��4�Ūl�a�6̤�;��F��ԧP��#�t��?����{'W�lD@� 	@^���+cU�caϷ�� ��K�BBX䀨���> ��h��7>M�6@�ܧ�N!���x�:� 0L��\��a1�ﯠɝ/6
�����0Z�H�x��_��]0행])!�3�Z��/B�r�5���JhD�E��,P�����%����ޓ�(� �/_��^��0e+��ب�]�toO�Z^�e�<�E���=n?��U|��.��2�t������h(�_�L�2x1'Ŭ�p��pyGEc��;#jD�X�ni�!p��O[g���ѱgAcʻ�����$��y���	xP=)�� V��&
�+R�vX�R��������suptͨ��H/c:�"����~ң�Fta�Ŵ��_g�< �J�: �]�*_�����q&C9���*��q��d���yi����T@����BM[^��>���ڲ#̈́� �������c�?^h��H�������z��
[���>d`��Y ��I�/�"ע�ܯ#����	Cl|ܺ�)j!� ]
��*�&|���(W�[��J���b���o|����[J�����o�-����t{ve��(����Vr%\:�q��K$��6ҍ$�6}˪Z��m��E��i'^��ןO3u�k�K�E��	bk�^p��p9�.K\,�=D����B�D�3�� }�.�����w�L�a��A@���*�"lN@�����#� � �}�M%89��� �*Ŗl����RPk>7d�Ҏ�Ig̱V�[1�0�9M�29�� �%rE���_�����i$�.�*z2��qG��{�d:C-���Ǜh�c,��*n��ҋd�[2�`�f��oIg�6=g��Yf�n�%�>x84MYa!"����&�\��}
 ����&	�E�X�C����{�h9PO؜����K�#�%�س �ٱ@��`q�49��.Y��fꔮu.�]vFe�r&w3��)��G�i�;�q�e;a��'�4�u��%Scs�ZW�'�c���}�vp�aw��RK�Z��\��&NVO�i��,c� N���# kxv�v(�G�S�F-*4ݹ���ޠg���܆6�<݋�i�sq����TZ-%}����*�13 0�)�qQU����e�qm�).�;���~_�;8v���bRUr@`��Og��SZF�}}	�&M�z���lR��};���.�����3�����z���uv���KT˫D��B��͆+l�)�-��L�Z�9L�ߌ7��r�.��o�W�P������7�x"�;g��sj�C5�W�e7�¯{��"b�k�,} ��w�gh�>��L�Ig)O�Џ9��7�ŀ�E)�{������i�j[��ko�Fa��[>��e���P�D�QQ4md��h���Ŗ-�in��=��3���2��W�+�i�!�q�p��q��4��j�n�^aEMk�k�x�ϲ�-�L�;H�uD�^��J�Q ��VH�R�.(�cȍ��ʛ�q;;c�ނIUn�xL����k.��4��Aޝ��,���Ҋ�^�nM����5Qx�.���,�'�9��n\�3a����o�Ou��bg���H߱�P=�bWE�.�{�P�����Tq(�lV`���'�]�$