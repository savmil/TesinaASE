XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|��"$�����Κ�D�d��G����q��E��r���TW�۱��Ҧԑ(A�_ձk�U�l �מGf =rކ�l�PPbDO���F�]�����@�q�'Z�L����D{�a�#��ݏ�B��D��y��A����#����F��'Qc�����lFV���Sb���ϧ��W��n.���Xty'eF��������E�K��+��c8ӆ�=�1�D�&7�˓�t
��X݀j0�����MC6`a�V�}I��� W#_��� Zq�崍��׾M��ޠ���_d��єÔ3ހ15��#�N�0�K���ܑ>����^��?-6{��_�Jd�`�Z�V��0��H8j�՟�����>�^�4SG��/���:oΧ���]��3��Qt%P�6u��!�y��װz��Zָ����4?T:g��w?sAΟ�X(��|���&�7�%]j�~G�`r�V;�����b��r��,�^a�np����0����ӻ $���R���T�.9��s3Օ�:?�,ׂ�B�|�0cXHSa-�OE� �w߮TJ�ϴ3��T)`쏍��|W-R�Ե��y��vŷ��e\�U(
���ywx�	�%�#w��Df�6A�C��m�Ыo>����-	���0]D�G6��+}���U�1�>�Pps��g�P����e9�r=J���]#J��d��ɹ���h*U���1��\�tG�OI]�C���.�f���~�J���y�L�b9ZIRV������'KR�XlxVHYEB    1602     7a06�n��<�5�w
ɐf�2N��rR�f/b��
��gQ��Luʢ���m�f7$��ę�3Q�T�C3�8��J��YkxZ�Ĵ��"޹�S������8�u�I��[�RdF�/���
�&��X��ta�{���aD���Z�v	�\�E�f�Vq����s)e��$/�C�@'�����7��Q`j�}y�&�Ğ��	&���!p�g쟊D�1~ǷҾ_	M7t׋�Z��=�&7���h@@@!�G�Qn1v��/��=��@�M~Â�cv�5��ۑ�T�'�7Ų��ôi:E���B|����� P����Q���.ci1+�ϯ�,�ު���f�.8t[=���8[�i~�l#=�-��Q�1����%]Κ~�1�{*�l9��ԣ�E��X�<O�Ed��{���L��6����c.�m)�P�(|ӊ��h�i �8v����1/����-x�'>��%6��k�/%x��Ȼ#`�'�� IFFnA,��弡�o�	:9�s����ʍ��<.�d8�`��Ϟh�]U�q�� ���@"�+4�I&��d��f&H��A�0>͆���"�m�6S�\fa*�%�l�c ��5fU�BLk��p��V��#��m��v�Ҽ��q�v5� �˦jo�+u�1������dҞ���[����B5�YS:2�^��%�Ա����:�h�kF���R��Q�o=CAZs�zw���4�ݴ��$_�K��:'�H2��H�~J4uG�i|�gz;^��9+(��8mע�M��|٨�Y����.�&'�na�>�J*w��>^��@��[C�.�lu������u]Zm�a��V��WM��^g�,�3�}~=���$�sBM����Y����J�=��^\���ӎq��T>��5+ �rL�(Mu8;<���RB��`��c�3�Q)ǲ�H�������e��Y�dN��J̄�<ۏ�U'&;�tmf�Iv�����7m:��(/a�P��?.�~eI�=/�_2%-����ye�>�.��ܨKz ��8���yj�=i�R�VPUɈK��ɾ��K&������%I����~D���"|�;��<�h����Q=�3�l<��(�&�߾$���ac������]�D�u���#`Ѝ2r��r=�\(������X�+���Q�#;�Ú#��˓.��Te�D��������ͻ�x-��C�]ڎͷ@�Z4/�%e��N^��ɮ�ޯ��J��mrJ7^��TW�HG��a��"���֪�D��7x��8�:��b�^eNӊNoN�(w9�W..Gi�8a�w�|�1��W/]�bQ�4������g�p$�std�H	��䗍�[�!H���b_�t���%p��Q�ˏ�zQ��Q�@(�{�w����8�d6��7�-jj���~��ز*�{W�"Rg�B]hl_�Vu]jF�_|�Tw���0G�.�@k�k��{J�K�����ΥG8*�]q��jT�5���y�Ri8����rwK��JB6f���
����Ƴ�w�~�D~y?(X���Wo��9�YO�X44��t4Z�u����x@���Z|Z�*d����C����Ǹ�L�ު䦫S�b�e�t�?6/5����^:��nJJ�?a0]"A��x';��с��.��t,��Yd�ee�Wh��O,o�����QfB&哣&B����)F��ǵ��=+�"*�;�jhk�٨�H�,�H�`����U�i���Y\ �&c
8��iY�J�}�"6@����w�dq��`G#���Kg����7�v����bs���ߐ�(<��:;�u4v���̏�B1v�2Ҩ<� <�-�����6��q�jf�6��0d3~��?L���_�#`��}G�}�_,�{���X����S���ܤ�Ig�T�e��(&wV|js��>7 M�i`��bDX/