XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^�@ڴޛ�l��֏��)��*7��o�%LAu�[�d��y�#�L�&R���%KnQq��q�Eq�����˃ڔ�z8����i�U��gl\`�]�2̭�����U#S�G���To�� �m����IK�Dx�Ɏ�čs�D�]���� �� ����䴝���pq���ܦ��9�1�\8m��Zp�����§�O�*�������\L��֟���uC`����cuuӇ2�S�\B��D�U�|lr~��</�T+>��M��J�Q�j&��kh���~�f��N͕�e�`�}~߫
c5nS ������=��W�s��c:-$��dO1���O��^�T<r�G;�	s������n�!��ѯ��q�HI�ݧ
�g4�2�4 ,��8hI�.�-�����W����ĺ^.R ��?<`���g���'��(fMݽ�t�H�IM��d�jCK����kO���6�?�����`��QL�۴�j�Ǎ%�x/8�j��({�*i��I�g$K�m�d��
��;vM�.Y����o�;�L'B׳h�mud��X/7���0i��`��ˡ^߷+��EX+*N����k2�5m�m\��]����d2-AMT8��7����$��c:���l�,���tYMe7�8i��")W�{JT]�n�L���/�q�۾#�x�I�܎(xMB���_�'У^j�lܑB�o���	�L�V߰��i�o�9�zd�4wi�R�V=;���,�XlxVHYEB    3d5b    11c0�����]�+��7��2H| W���O��BA�ꁍ���ƞ
 ��nEK��0=�G�B�
�]�C?]�W���tq��c��!��R�(寓��~�4�fd��^i#hA�+���%Ђ��.�V�]Ij?~���ɐ4������	�1�u���^}�{�~&�g��^�"�����r��u��t#�8��#v�:�չ�W�_�H�6�)f�:� &��V��F$��/��q��AX;,5����_���!�+1�ܪ����r����ٞ��r����^t���E��-��f똂H';�tSc��Prh9U&��{
�Aj�l�t�j�"��|&2~�+�LX�&r�%<ڡ�J9`pzJ��xT��q!ZB��]��َ�rǊ\u��M��<����nh�(_Q��k�h����j�nr�|D�CO�u���hV�1P�����J������g�XƎF����ɼ�*���k���7�� ɨ�72|�{O�����fZi�4R��6�E^�4:�W��+��t�HX�����`�!�����4��8N��$�+��[�~��3��a/~�{z!3�6T6S�<��sK㜠�$Q�W��6�����!��p�?��|��d6�s%8�a��њ�͘���?��ɻF����� s�*4+�,�h7�'#�Kl�y�I�HT(�5�ˑ;��1��S�����	t��b��R&3v�H�^��4�^�V!�@ɫ��zۤ���'/�S2���������j�eIj`����R9��>�M���2�	��֯�n���E>\ [��|Q�I4��X?��@�}�=����U��l/Ll
S�nQ���ҡ���qX^��uLh�g�$'�T���=���i���� �J�DV,|I��Xo`I�4��a>�O��m:�B�`a%h��nf�7?8e�"���sUEV�1s�(�Mo_q��Ɵ�Dj�p��M�;m~�Ȳ1/�:ÃF��=R���d%�m\C�+O����Y0������&P�Y��ގ�β��:n�%+	�e
��a2��sr#����O>;�K����=u�x��I6Jr�ڿ@0�� RW�Z���*�ݱe��j�J-J�O��:c[n����$�j�sp�E�]k@	�n+����Y�q%���Y��	1�u�����y��k�^t&Y/$u�Ф<W�H��G��v���T�]�D�j�`�!�>���V�^D	�)�U�:�H�Eq��#�\��7)�T�7=�N����
Z!�3�^-%�o�������A��vk+�a���2RR��7y6\L�e#�����o2u���:+m
5�w���P��'^.�`bƚ(&}ꐺͰ= �����r�s�txP�e�����20��;>}8�3Ԓ+�c��V��ڠ�$�ڑ�\!$������Ufb�,�g��}�;�8,׼��tš��8�6�`�w��	�U�ww���w{0K�[#���z�'+G��2���� ��_�|?���dN_�t�d�)K�OZ��K0χ�V�ܘ{��Ҋ��aP�C�,��d�� �t��B�D�9�Y�8����� �7��$肳)߂V�4���X'�w����ɬ�I�"'}�K�-�۳��5���vY�` ��%D}�4n#nkO��1
dC�/��f۾L�b�	��.
���y�d��e<Y/@���"��VI3���~}��n�蔆�S����n����3�,�#fKA����-t�_G .:XV�$~�w/�M)֒4f�+��^�J�JCDh�ځ�@{{ySm&Nr�2����{e�fci@�O��*(����L��t��%�k�RěU��-�1յ�VӶ�O>?�����:c4l%���J ��e[�� .�~bҠ������҈����gi5�
a�]+�g� M+�B��j���`�XGp���*A��w6�pEq�x������ڳ�"�-��p�L�c����)I��.��<�*�R�UEY���Pϣ����K����%/�B�.�-��	�F�D2'ō3�N�R�_���+�*�h�7m��Ա���v����q.Y�^��?��#:�(20��Xz��|���F���6*�~�L���,;��0��u+�`6d(a��u�C�#iA\�`@ڍ"�������,v	,;�fE�xw��,� {0��(V�2�������
��\��KW�2�#L�Wq���s��Y&K�")�sw�p�����a���x|;ȕ��,adĢX �
r9-�>�A��Ȏ=?����N�1/�m-���h��<י�g�m��ރ�'�i���$�k�M�.����(�,�}�+�>	^춤'��'�i���o����4W���R��Fpr���i�8�?E)/�gq���G ts(@�R�慤�]�A��!u�~w�乘
6���7�4������y̤��a�6�aЌ��C�vOwFh��w��+�p�P�A�_ ��{����=X�N���<:`����ki�O�d�a�N�q"�K�04"����xZ�Ge&M�&��	(O	+�;!/�wbw{N�G΂n5/��! ��������ܾJ�5�:J��ة)c<̌Ny�s�+�<���_�ǹͪ�R�Jth�3$�P�_I�\���֊q��N Zn�=өa<(W�F"�����Lp�t����s����S=�a���EȾ�k���e����A�\NVk?pz(��#�L^����s��3>�X��|�J��m�IK��y�ҥn�}P%D$:Li�w�!�J�S�o�{
C�{67H���-����5�t+� �u�ѷ�i䧙��3O�b�Q�WYx��::@�]���~欄 !msg�����o�`�e��
"����tA�Q��W(����R�T�h4+���b�
��>����4�� $�r���K�7�����)�T��#(�~��J=�s���g�Y)M��p�%=qK+9�a�4�b�g������]�Q����@��\�i�^Qh�"�qnZ���ak�aw��YJ�A���3ҧsU��E��?�O��8zL	��̮ͯ����eh��N�_�Ī��� >c�Dq�ƉD�x	3��R�s�0ug�9kb�0 � �9p&j��.�׷(�< oM�r���o�D���x���y��Z'���ւ��UU���M.r�T�	�M���Z���D�����mk:ei��	�|�#�ݫ�f� 't���]i�8R��=`A;Z����ߚ��2˸�jY�~U��AJ ���ެ�9���y%!�F�i[I�4x,�2������#o�pz�z�i�u�$~Do���J~
���م�����Z�
{s|�Xڻ/执�ާ��(�H��k�y�xE����}}z��ec�qͭƝ�n_�{O�wk�'�2o���X��Ʋ��:{�+C�&I�������l�LAb��n�'d��1!Ts���s���<�I����t-`�w3�"+-B2�܂���v�ġ�<�� �  �D-)��I�-P��w]��zӏz#�i,��W�W3�V�J��@$�����Cm��!� �Jt��JR���i��?�+�Z �$7'V�RjB8��p��A�/t�����1F���ǃz��2G�w���BG�0?D(��>b�[D�8���	5E˳���E�* CW�G�(o���O��/�$MOX�)v��7R�Qy,B��}G�_��� �		3��Fĥ�_ԅ2��zJfz�N'b�׀T�?�a�����x��Ta�x�L��-*�������zK�,���Cׯ�҄ąnsa�
ŗ^��/Μ�)ASYc5��B�(�A�Y�0N7�qmd<�XC�1�X���yWD�3�����H�U��L����ٚѻ���}���y?t	�+4�(��nQ�ڮ���k��񯦳����x5��	�I����@Cn��	�}��m�( ƹfb�"�)HTjm�Ô+֔�+Բ �Ug#Pu�:�A�@��j$�G�'�RЭ��fT��uz�;�I�@��� L�8}�ǭ��O2����vбD:g�L�Vx.��P��g�@�m
�/
��<��>���	z�ԙc�Y����~kM��i�2Y���r���l�k�w�w���Y
�J�t0���Zjy<m��W�����+6r���P���_���FK~?cI����J�c���t}��1�|�¶�Yʆ�<��}�'���S�[תM��>P��u�Qޠ��Υ}δ�iZ0G�����|C����:����ѬH*44ɴ9���c=�9��j^T�=! LR��TȧK۴� 0K�:{�Q= �N�JH�|���t�~)�t��֓ډ���.H�@�9͕�v�]�2�G֌��fҵ�	(T�`�E��qj ��Y.ӳ�8��,���8I� ��)�����~C=^¢��%lp�� )������0�
k �]=�J?�\,䩶L%=i�t٢�IZ����S���N>��mM�O$i�\40xXL @򠵐DO��x;
[N��u~�yr�