XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��҆t�4��Y'�/Zo}q�e��H�f���I��g<�^u�����������+ ���sp�*{����[��7E�R�@gW �����lD�.H�W�{ay/+D�!�.�F?����\4qg�P�bd��"5���f�$޳�#	9=3�Њ�A�x]��C
�?�8��)gX�L�/mE2��:��\t�<���;��	T'؜p��s�F��娚a�r�g��Vټ
�+���+ղ!��"�D�"	�6�GMo6��>7�MoHY/���R�x�ԟ�2�2��4b}[}��o�xk�����rj���N�=�����3ڇ�h�)�8m���x�]_���8a�T�d��0�<<����_�@�ޓ*-
������BǞtcʖ��	͸�q���	�i�p�	��p��eq �e�DOhl��UP�G5�=z����r*�w���ph(��ߊ��d�P�2�I#a6$S��J��)8��{�$� �(}MK�����%�2 �����M.�R�I?�h �v�/�C��SD��pq/?[Z���TY�M̺�%0���7�w]+[���ܘ���U��_�x��`D#�ܓ��V�'�g��� �8P"��\�ƜQ�����2�f*��u������?��_w>B��*M���M0��25w%��6�Q;�2 ��21��/�#�g[���2��*�͑�|�A0&)���86��e!���3jx�M����mX�T�������;���ֵ&�A�v�	EXlxVHYEB    6e28    1620�����K^NkMv����#�h��\�1O��H	�G�z�+�
�>،��^�$�Q�����aʛ!�F�p5<U��"6)kΜI����(���jI�2��?�R��|��(��Z�Z�q�����y�x�t��3�ᇾ�xy�j܋Y�*�����m��_�'���;QW�����U��ui4��{�@��j����c�D�W��c��^:`pÆ%��i'�!ٚ ��P!�~*�k:򣩳��-�մg%��o���p�;��]�\Î�����J{�/���m�H���hu����'KZ�I�X0܈S�n�>sy�3'g' ~��|� 񉙗���ґpLr�&L�3I
Ė~:F���]�sw6ɉ	�O�@�� o�P�߯�OJ��**E|.yO��Z�-_btV7,�n�9o~2��N�ck�iN�>ŝ��x䟶�������1���=��~� �zܷe ��LF�}�����[��[�<=��i��[3�i.K~�2-�G����x��pm^�Ֆ,W<܎������Bl3�2C����y��;K`�d��Ѭ�Rxn]�������|o?�y҈ٜ�f%��L��֮QdϜ��C�=QM1V����iw���y�	�"�2���@�-�¿|@���$�G��(N��'���U;�ܤ�^D��PE�?Fh)5�}!�`DBĊ��s��C��⑛L�M֧</�H��Y![��E�|+������Qd]��ά�����߯y���ù�`�!u�K�研���	����sەV�0˘�t�Xu>C���)A�0�P�7�;
*iP�	,���q��tkb3�G8���fǾ ��L�t�N�Yz!;��3����'�x�t��_�Q�W�Fڶx�)�q+nzA�%?��:�ʯ����O��NP�|���G�`�4�D��h��8��zb���:cv�QBѕ*���S��JLS35F�,;7�GV�.���1�}�-`��[A�U]�i��$�qB��$)���Z ʙ�"θ�+�B�V=Z��� �%���U/�T�����wŎ
Tu��I4��v��`'x��v'��K
 �Lu��#��飑F���k�LQ'�lȓ��N6�g�#r;�W�2~W��ɰ���?��m����ŏ�{�4W�����!� 6w%C��֊㭪���ˁ��=mW;)2,����T��84`��W[Ҡ���?=h�hM"�˘���3������%�ѫ�m8G��۲+y}e	�k �V��l_NQ���"o� �J�g'��w4��<R�?r� ڌ�q��6�(���Zj=����;j�W��?(m%M���� t5y�����¨�M���g��ۚ��N4J�p>$�^��>�f?����S�w
c�6�Ǣ�5f�����xܝ�گmmF�.������ėW�9�td�0X�qW�C��JOv<�geX�_�6Y���QH�v�L�|Ki����Ti�f@�myU�N��SZ� �ۻ"=�z6��?���>�yz�&fh���3|r2����yY^{zI	��_�sK�&��"�ǌ�7&*��AM��Hy�b���6��Ѽ; 	��I��z�zJ@��V��ܣV`*�:��d��Z��~��F������k1X�~F�jF3ۘ�r��*�hlc�ǁ���c.p?���<Q�'����	�=M��;S�w��V�-�@E��E����z� U;�����Ә/]?v���뙀1��4=��B�Q-4��B��d�{�v�Ɉ#�����^B�ɯǽ�[h&�$���d%����-���jd�B�*�Կ�2Լ1?r��-�)��,ݮ��n�Id~��՘��ྫྷ�V�v�m�K��@:�(�=?�X	ס�o���ct�:RW��'�Y�5�K���WR��ɇ}���W!��!���
�gX�\�q7����G��L�7*5��\��q�B��,��1"X&�Q@�u��3�KИ��%�ݨ+�p�s8&�<�� �a��/����\�j�D�/
	�=�/�q̏(y?u�`���@��qsHτX7�!�J�>[%�Ss��A�(�{��90�Ù.�>@�f���̚u��2@�%Zh�?����Z�+aN�y��l��Y����Q%H҂Fm��-_�������RJf��y��Ҝ:|�{����D4L"5yVW����ܳ���f�.�Ҧ�D�0�����Ù�<=z��n_�Wd ��{Cn��@lS�`7A+�s�6,("���'��Ҋ%u��WЛ�'�I*^@���/�K`7�]�ք���lez=<�� �o���܂o����s�8�Z��9�.����d�]��BBG��b
����t�Ikc�w��G��X#��)��:PG��>�c���[����8�~�kGF���QݣE:�>���+���!�ȡ�:G4�����`�"��WS�Z���l|Kc�7�Φ:W�E[sJڶ>|��l��7W�R���q��k-�����m�:�h��	�h��%�h��W���I�f%^T�x��Eg4�c�b�'�T=�ű���+��0�k�:Q	�n}���ݏ�"�{������(Y����!I�`ǝ-�۸��9���32�
7Q��Ȕ�'3�2Y?��7��� �TE:v�����Ç��Y-�@���L��"'9a���2k����j�D�W�D�pU�|W֭��RF��y[&��|UC�ܾ�f#�''������)�2ܻ��d]J
�&&ro(9�4<��W
T�'L��|6�51�B�z�dbD�q0,*�`HH�����PU�� �������E�����˱GQ���#!J5�ڀ���M����;�[�����$K�iM#�C}�v!K�?��+�^���!¼��N���A��E�����Q�_��5�pp�eW"F_\o�-����g+I�ޖJ=�Zέ���Q+ *�"���>��d(	-&'�P~�I�g���=�����	��S��/Kh��(�G��T��� �f����M� ����͆�)���tJ��P��$,d-��پ� �Y��_PWE��g�o`�I���g-����Y8fl	H\���`�PU����~-r�/'��3�/��5i#�Uެ�2�k�ϭM���6�eּ]Q���i&H��&���][�'hA10�=E�a��Q�Ap#�oD��(	?|��gO��;,�8��P3�,5���T����su�H��VV����wx��SZD�O掜���Au�����[2I�e (��u4��ݗ]���s���8������ER��I`�� ��~��G��8�&vg6R�DDDF���;��D���FNo+ۈ���������OPe�T_�7�W���r����T��[��4�}��9�s��%6SF��J�C�;~B�wG�U�`���3�|��Ø�o �6��No�m�Q鎊Ǜ��X֐��޵�Q506"��I͖�	/�9�ݵ��9��\����i�f�W�q�vr\���5��L(�}�ٰ)��{�����5�E�Y8w�������ti,2��TcB:����Su4��ǋ�����o��/���)���j���ٖN"����ѭ�)_�a�!q�����6����Tb�\:3�`6}>>�@�k���`��w��㨚:��M��e���M�&��d%r͢H�3��?���)��1��K:��� ��`j��l�c�JW7̓
V㟒y{�V�ֆPw���ú=���E��S�` �]שr4e��{���Ob*0m f<��P,�q��6�3��ƱZ�Ǘ�����X!8G��m�~9,���bjUш�	��lٝ�`o�Tp�7��t�#���%���=c��	�&�R��h�b:8��^E�9r�/b&2�_������ypRZA'����c��\m
� �����@m���.n9Ӵ�+����y��v�N)8��][wa�9��"���c�0�Ku�0A�����	6D�"��(�+��y������� ��u�D��I;�>�\�EXz���G�ݮ��/�@@f�&M�O������ �3���` ����s� �̩�Ѡ��W�G��_�^��El�m�x����K�0F� ���Y_����&ck��㌬��V+�]0�3��Cޙ� ���v��ڮ����WH�u?!�ƭQF6h��ۻO�
ۘ)�W{o��_��8ڹC�fP��������z��XL���e��,Y�� !E�MI�� �A;t��j!��3��r�O��2�-�%L�pEU��,��n]-��TI	"4\�nP�.�0N*���=�2�pbC���H|8Qb.$�ٱ$�I�&^��+w�/��x�;�V{^�!u:	�?�^`h���;N�� 6�(<�����Cެ���R�>c�d�4�D�!�d.9�3w1���=i@l�|�����������O\I� x`d/m�I*����ɹ����[��L��ca��}�'���-�f@#E�*,/����HkӵS��Ή�Xe�!�=;�C��煲��y��TB������$��k˽o��t/��P�;�E�
S�<�Ys�F�����/���?:�]R�j}[�ۤ��� ��Ş�� ��wT~7W0�kK��:�L���z$t����Nqf�>ybS�Z�.�t�~�ͱ�ې��4\s�C�_Bb�(��&S��x�(9�T1�Ƶ�V�Q�R��JƢ�6�U�Y|w\�&}Y�z)N��ۉ?��!~%�+�Җ�2��gZCJ�2+�������'���{oBO��5'��14�����!ԧ�V1p#wO\�~�WRba_;u]�(��D�� �+P64��S�4��(PU���e�NQ�M9	(5�u>H�B�*�0���S�����j"������n�|��-�"�="�^���o�����8�V=�̉|M���������V(�j�ЂoI]X�'A�L+����W.�O:����%;$����&!�H&��K�GD���aQ���"v5H�k2�W�G3�:�e��[��$D��b�DzMA�x�e���"�?�;/�ܘ�(lƈw|�ސΆ���nb&x��ݍ��ɋ�/KD	9�	<|j��+���y���=�%Ri����n�;�Zs�1�O��?F�(0�zYb��Έ���tZ�5�(B�lH\���[M�Z iμF/���y����k)�Q]��}T�o�{M���9�#*�r+y��hF�|V⺈�����0�t�E���Qσq����0L /�U4ju��M����쫩-C�s(�����8���M-x86���_�B�)���Ԭ���Z _��=]���Ciw`���:����K����G��%O�]��9��\2J�}g[(�z�X�C��<�P_TG�f���Xα%������Z֥��� �_�]���n�8��;a�Q��)�����J�>s��.�BR��AL���%/P��HO�j�De�|�E�i� �<}��^��2��BI/�[!��������͔�R`ٸ�h�FI�{q�.��@�h$�9T�ҿ���ia܋�D{�#ܛ4����ќU�@�* �	��{�{�Hq�;���q�e���w?�V*|X�ӻ���^�V]�No<�� ��