XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��vD���j��J�Ю��.�<�#8gL��D���^���A�bE\�C2R��3T_�3�)R=�̂��ОAv[�f�p�ܒ�F�J���%���ssuq��+�Z눦�����l{�b�?yru]ը|��c�����c����zu�%/�Oϣg߫^-�.�Q^���K����Ixn�H�P��,��w��ꆱ�H,
B#-�Z$�����_�?�ʫ:54�!X��`�����Ao��H�^��a��r�Z�;[G�Eۚ�U����1�X�Ǣ���ܢ�|�8M
���P��Ai���Z� u�F;��܅�'�4��}?s͍���7�p|�I�R��̐�/>E���֋�9M�gy�߆�>���]Ym�f�q3��0raG|�G<"��H��}0B����
"T����.3�.�' g0�9��&o��n�)i����rk)Z
�'i+��C��՝sS�C�h(�E�é׸����:ܮu��yϧ��"6j��j7%G��y_t�i>Gm3$�E� ��<,JHp5���o�y��]��QȂ&1�8��6A��i��jA[b�|���EU�D=CH%�g�����Q�[����}ᝄ
�b&گ��O,f��], A����!N�u��l�����#�@�l�����!{��?;?.p��#�Ÿga׌oUH���0�����'b�T�v4��땎ٳ89�ts�(����4��_濡k����tͲAu�	�+K2�η����B��TR8��C4*��XlxVHYEB    5e75    1150�Jd%�z�S��!�VQ�2&�5���(����N+ ����"8ž����^g�`D���8�Hв���'�Ԇ�"���`%���&�^����6��ʇp=�bh4�YC�7� ����ċ�ߋ( �[锝^��hG�*�����sP	��
+�Nb9*�e)tTcT��%�4���Q��[w� *����c�|:���~i�8��U����W�k�d�����b~ѥ|u�[5���c׀�fvg0�*� �s��ƥoW<�.V��i��\Ԃ�7I�:d��F��H@X�O�f�@4�SNC��ͨ�<��O�2��1�F�EI��Vj�g	s�z��t������&�K_�E m��Y保����;ٛ�W~uv���769�M�+�~I��7�bC����<b���z�u��[\Ŕ"u����Wx(I>$W�#���>���W���W5�<�Պr�p��D��e�h����F=�a�{x�K3[~k��Ÿ��Tܝ\������*�~�OZ k�S8�	�0��m�t��.5Z�	�G/VVl�q]�c@��i���4����]�=�$��#�W�0bZ���{�zL?��߮7�Q�Ӷ%
!-�0Q$�~r�ݱ�D��	~|#t�=m��=���C��[o1��(40mf�imK�f|����{���׫Db�K=��k	��\�շ��(U�19 ��fN��O��$�hÙ(��9�EU��+kDG베F���9'&�t��4�
���u���o�]�&��&J�ES�Y�*���+[~1����P��(�v%)�C���']�T%
V�S�cuLC�S��9�_�.��(B��
�X��L��D�圑o$u��- ���{T�e��c'�^���)��P�w���������(��^���^�:�IMC2#�x湱y����#�2?(�i\���!_蒞s����^F;dYoTG��K%��I��.+��NתK���uܨC�O��d�u����uxh5n4��y_��#�9�7�mbGe��]:�Ni�F�VF��F����)�)U�}�l�2����h#�y�ŉ�?|V��m���
��4�k��Us�~�;��4
|�]�oo��vֈ�-˽�f)��o����-D����
���ri�qؿ�(�Y�Y�t6Usʏ�%��������g	?NJj8nw�#�j{g�e87�JOk;<Z��)#;���Ĳ!?�m����~!�"�V�~�	�����!��|~E>�cAq)e�6�t���(P[�����!�G�S��F�\�����h�C��yp���*@aM�>A���e�"(����,a��]$�mr�O1?�����w��\��I?f���O�ސђ�� �c�rzpD>�2�@E��?
�X��#L��E�H�3��9�>ߧ�yB��m)�C\4����B���A�pS�l^�����:U�q��&�,r g��h�'}���|�:-��z0���_��K���>z:|�:-Aa��F�1���rk	��� ~���2)�]wǐ�&s����;�����"h	;�D(8|�6O�L�ڜ�n����o��Y@,����Z��f�k����oJ�F��F4;���#��4�q�v���2,��F'A�07n�&Ll@��X9��,�b�xe 㯕8�vEɽ��lk<B�� �.�S���I�
8x9�r��ߌvq�kȅ�$XO���"�dZ�65	{}���4��#�w��I��BT�X+����;�7����m1_��h�'��_�a����)��}�Msb{e���1����8���+�iM�	%��>8��f�W%e%��B��+C���o�*1�<������ʸ� ��y�tS���e�6�T���O�h��!p��P�na�;����o#�E��>���E����Y��-�ȵ�H����SǄ�%UB��/ � ���U�w�1h ;��F�J��n�G����>F��E�7�C��ҋi���(�'�p�̡* R��:ۍ �0*.³�ƻ�����j�˟���CB��4��(���i�O��ޥ��_ٳ��qG�a�^6c�� �N���?8��.��pt�1rZ��V�[��%_K�r���e��lO;�x&��F]�Y�>�mK�N���Mܼ�}Kƿk (ܳc(]�[a��<A�%T��I����o��*#Z���)��#K U��\ɁB���+(����*�n����2�w2Wj��}@n��V���̳��z���n��!�DrA�[޷.�=K�߰���
d~����n���e�5�y������M����,-"�9��I}�� �-n��iV��Eǽ_=�u�n#I�Zxh����X
�"����?��_��]�[�9���U�{�K�ъ�,�$��4��z��P�͊�	5C_�!cE"#��B�؁��d흘*V�Jn��}X����*I�v<���\�����ŽV��'��~үh�{a���k%�O�\�7K����i�������t��#A �_*��8h�	h�1t�x{;���.���i޼u�y�i8ڥ��)�@b�C��u���E��u�����H·ǁ�������a�Ʌ�e����jfP
S��H�/y2�q�l���6�v��=`��N��u�l��Ёn�YC����s&p8Z��@/�аɨ���uk�^?�=��%�Y�X�Y�;N�-��[G�Lf�鵶Y�-$E0a��y�ނ�GA��e�@��;���Ma-���pG�S)ĺJ�,I��mj �?�4� ����G�x��p?e�H`�TF����*.'KQ��!��>�S^��9_�J��� O�����/�s��@�����j���s��{l�����]�l���� �[��cU+��U�XwNSeZ<�{��L��J�r�x�*1���f����̛ħ&���[x�O�7��/�5XN��]�~�ى����m@�W���wO�)i���SP�܍^5*�pД����y�{�|�S��d҄��̮�2P�E]U�`�L������UTO(���N��f��+x�5���n���ʚ�޸-��#dS��9)��7��W��8^��B�D�BS�Z�0��KW����+x,>�����^k�-�Lp.�+�Z�xh�����$
-5�����}�,ȐW�(}k�Kxw�������o�����ak�RG�s,�������)�"�ޮ6���c#<C�g_&���Z�ng�������u���NZ�&��i��6<d��G�x�q�􀏖�dp�m��W)��tخo��VbU⮿�;Ye���ER��!&�1���.5-��$p��#,
MG@c3���Y��N�8��^,�EŚ��f/͈��fʯ�����g~���aBi[2����3�J77
�	W��LJ�)k��_���r$�S\`ˤ&����0'��j��8:�^d���̧>V�]�t������YZWI�Ӳ�^����=���C��v�	��ۢ��B���{��ع���.F~f``������B�-�|�����m� m��o����%��JC��Q��
�k���.���p����tgw�y�Y�z]y ���ss����ͫ2�Q�E��x�O��K����׼�k�j@��Lc��yp�������1��}+8�K��MR�����*�L[i���R0��Ԗ����X�[ӂ�>���:-�,�|���>k)��LL�En���*d�����G�0S�9;͖	8\��yK/n?wE�s,p�c����V���GS�w�u�_�]�	]rJ�x�̀��q�L㛵a�>�+r�4��i�>|��
o���uK�{q�|�t�����Wy�X�2�%A�[�x�����6�m��8_]�rn�����oR�������4�`�q�����VҾѡ�8c��Ot/����zZ^+đ���lIc��t���rFƠ�[z���D�>j�>-�iL��f��E&���D��1���Lm�nd +�ܣ+o��a�B]&����kg�O ��6QSBX����9*���1h��0�eQ��9�t��dga��d+&az����������L]D����
|7ChR��O��/�O��݅P�)�_sʋ$���
;F�?Aß;����t?�_�;/�L]���]�wѴ\��s��s�Y�T�1@��K�|=X)=N�G��0����-�!�?j:w�=[/������y�-���4)	&9]�}oF���E�϶b�x"�2�ɗ{r�[Xw-ep����#�\�&�F��<��mE�ǲ��#!}8q㬇%?4lI*%�y$�-9���S�G��L��k]�'�ُ�k�*	6>s�H�)�W,U��[�u-_o�K8�1��!A`�� !��|��&�-�