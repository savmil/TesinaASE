XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����9H�d��<8����P�q^���v�Gt>��Eiw�%mJ5�p*� 	uGp[R�0ܢ5�e��|�e��drv�6�Ԡfq�,�X�8��qŝ����R&p�x7CQq0=8�4�ef��d��˹�$bUyM�(8�mrw?Q�V;��L*��(O-�yik�&~܇˙����a��L?������q�ML7O��OK;+4r�r$��;Ju���a
24}b�6�Hm����f�T�>7zS����ǉ6���T{=�38+�CII~&�0U�sG=+RU�ېE�:;0�*��OM��g�/��h0�	�'�3U����N���ʁ?�>�<g�z*���Z�.�M�S-���g�������1��^܊�*��e�[ȗ���Z9R�y|(��1&W��M01�ぽ�̑ȿ�oݙ����E��J`�dD80��Pr�y���$ZC�|�0�6ފ:z�d��(
����&�9�������Sz1<���.����	/S��6� ۛ3�ҝ��r���Q�����t���/	���n̪��h�>���;7l�L��5�7����v�3�v����z�J��U/�9���./B���[sN�����y�d���â�=ԫiR�����[�ޮ�� �I���pWW�����GW��pݓ������^�j�d7���\�sA�;� � j����&˞��wB��P�X�Cj=����������P�G�V�xNI'v��g��*ޕ��*Z�C6{:�����5?��$0v�M�G�XlxVHYEB    4013    1050��L:)��N��>��L�����'ùZ�3*7����L.ځ�jS�&7�b�J�Kdg��@c�ū���i��{�U�������q��D~��U�|�~r#���t���_6:~!YX�5��̻��ږ��˛�dp�����t��	 >�e"�ێ��FY�4����g��P}:c~�I^߬�}�E5J�e-2a�H����e��,��;e�0�r`޳G�7�o�ƞZ��H�?}!�V���7��T<Jڊ�:K�[�[N�"tO6d[����>��!s���*� �%'R�@m�#�I����f�n�Ek��Na���	�f�>���e��]�,2�j+n,ʧ��9[�$(/��j�t�z�ۆ�N6������Mt����M������t`���bZ��aݑjh"�@Ɵ�'����u�
��z�唫�`�k8��]�;s�V�ԡ��5&�V�?ʄ� �܂��aZ�'�x��sc��k ��9�A�B�
���QP{���Zx6�r��[ņN�✵�At]}V�&{17	��ѹ��5��ǳ�; ����j��|�����m:�b*��0�F�t���]��v�X�#֊��Ũ����E�~�
x�y���۔K��5�ClDD]����H^��(Ul� &_��V�MS�P�`v���m��2#��<\s��>�3?1��Zn��hGrkmeZ8J��	��*qFp]m2o
�U#�,*X�G�&�zo�d�-J~��8}�_����C}^uB�G_2�0��Qu�A����+�H�4 ~F���j�0OP2|$q�V�PJ!�G��]�ҹ��/�	�^����h>2�8�q�f�8p%Yh�L�H�{�$
$;R�k�Vd�k]��S�&q�IFP�-��y�Y�N��)��)"���Ӆ��z�>�~cp��fT\��;}�����kc����q��}P��"��Ee� aD(�>�P����Iil"��K�e������;d7�[<�H�=�dJ�JWtvr�	�伨��4��L��&�
,;�d\��H�yO|�ZX�K�n�������I$�r���Oe@�K)����?�U�e,݌4�,��F%���ވ)�����/�[�51�5���W�A��1k�_z�w�&���9�^Y /.U���T��z�08��1��^���!��I�U^L2�O�	`�����6�M͞�vo��YoN<^�?�$��y�>B�䨉�Чv@��X�^�]�{z�ވ��+��J�YvV��.�s�#y��D&|Yn�9���Z�t�j?��N���0OE�W�&G����|`S�0Meo{�r��@�$�PV7Q_�� K	��e�q�e���Id��&^�]��MP�no��k�O�4
�c�(ˍ�`a�u,?�1�?��ː�i�_�Ob.j��"A2X��	e���)LY<�ʆ�����o���kLHO�A{���:�1'�S}٣3�_������@�+��:��ĩ1�_�A&R	"�$�Y�;��h��S\���Ě��a1�кSe���� �Ԙ T�����x�p�/O��3�#P���^�ԴA'Pe�T����m}h���S܃M&$3=�=Z���͛Vű�����D]���4��Vx��C�E�
�nY(�0[�l��-�NXlmw����;8������]l�0�J��V|kd�R�ؽKC�mݷ��bd��g��NzR "�!1�i�sd�,�>7���> Ǌ��\����Xt�t[I jЀX5trP��/]��d�3w��.=��7�ݨ�iDs�"q�z�
������T����\��!˵rW�%zm�N���j�pnk�1
��}�6�����َ Vh���\��9_��u3�P<ez���	�]�^� O�� �g��Z�#��Lk�0/AO�U�v�nһ�@���bwwNyJ?���kr�6�~3$���Σҵ� 3�;���q:���!��7�'����w������$1�6GߪI������n3����U��vȶ�k��pe�������;�ֆ4(�Vb����程���M&�=��&Pn�`��h�i��_������s����6��"��>u%[�w��e���&D\�.q�i�U��@�5�ݖ�`��>˲<
�ɵ�l�����ctz�4�wa8��-�p�C[�꽎�I#*�a�GxD���]=ϻ�{��p����uo8"�rd�@��?���E>�}��ef<��H�O� ��J�P{
D� d������W �߂���-4�92�+�lN^��n{$��9��`49hΣM�9�S����k��X;5�`r<��("Y'�ҹ4p�9Hw�s����}��x�lC!�F�y}'�)�b�����I������U���hώO�?�~�[רJ�&�����%�!phR�Թ#�|�6�H[@@{����C�Æd�\ۧ/8\Hm����l٨0!5�#ȝR�
G��f��H�O㋝1�B�( x ���[�p�V&�S��!:g�[�D!�n�c�yՖN5�&���T\���؍d�jYgX�Ђl>ӷ���E%�r��F'S֮3����̗���N�v�����h�3 /��#�����n3H�6��5������s��k� {�ՀJ���#	)����P��r?�r_6��w̨^��q(@}�!e6���O}�Ґ�w���"mV����wwtʄ0qz�MUMt�,1����z'���w��%w;���<��0;'���\9.(U����Y�C��0���^g) 
�U�����a�+�S	��⌧$��B���!��]P=,\a:��%�؝-� ��8	�������DT@j4wt����a��
+��Ϧ �p��W�o��E���A�����lg1��-���1�z[�iV*��h�/���L�����
�L����A�N��K��L��t|�BPz�
���|��h�`�kt��<�즺�"]������6���#�QHY�պB�9�{��=8�qU�w��'�T�3�JRT0�%�!S�=�;���./�]8�]>i�Q~�糎��3�~�x�.dm������;&�؇��y�3Tgk(u_�FT4>=�J��\���>a�q�=F"����Ir��T�>9�9�Ҹ�8��[)q�P1�{>�R4j<�{%�.[��&��e�[W�)�XN�\\��9��^a�h�W��u�}A�}q�__�}wo���A�����%��nUۇZ��w�����za�R�NKe�v����5S���A#�g%3h��{��	��������u��PU=(����\���`"sj�8!��2������s(�Çˤ��<+��8�X�B���c��%���W�>:��m\k�Rpw;&7�-�,��|�k�$s^��-IX��eMw��)���8
�o���#�ޅ?%���cf}�Tq�B����8�]�#g�$zj�Du��P�A�I��vB�W\�zD
��C�s���$�MP��P*���C��(8�b���S�֠��a5eQ��F�fg!��Ӂ�~I�߮���S�RH�k�u��/����W�4C-��|0����o)��
����4rT�(	`�m�̈́�ܑ(�F\[U
ĵ85Rɍ�Z$(Lw`kCaQ�%�����,/{t�
ݙ�e������DN���\�*]���AMC�%JT�Y�W�J�����Um���H���8	���R����?��m��d�b����k���3)�\.�TQAy��[�?���8)I�`Kh˱��q��gR;�"Wi�_� :�Tp��*���)�]�)=��$� ��3���%�b�W��j ���:��%��K���H��|$x�]���x��q('sx[��q�Bkj��vD�����rtk������i�'$8}�8m0� �	H�i�Q��B��/\:�K��E1��^��U�F�s?��o[N�:��C��	��8P���ƪ��j0$!O�K�D6E-�������׋'��.&/�����7��b���"�-v}�?�47����1�	m��S�0�z�ɰ�%�X̽+�L�E�U���4S���6�O�ß�c�$2���.ͭ�vM��ڄCq�|@�)��ZE��Զm