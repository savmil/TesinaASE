XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ݙ��I���M�{�Wh6�v��������Yu��"�n�|�&CWsϔ3V�2�"XΥ�9�U29l���Tm�DZ��d� $�b^��!�1�8�*B�ʺ���@��0��?��e�v]!�o]E��c?ʡ�1��.W��k��*jY�:3����W�����y,�t�ő�FM�C_{�>H��$Ï�2Dh�%�aa�(ɤ�_��A�.�&\p�-���i^��g(?�Ƙ�r�}�J>�Ğ�����9�@%/��QP>���e-u��<+~{.W�i�%Q\̠��J�����Ʉ4�f�xA�N@��U�0�a�
�SH.������-��))xu�~	��M���|�g�	R{k�m�]��!��N#C-���fv�*R���wqR^-�PJ3"|�a�����Ж)9�P�A��l�QIذ�|�$j��o~�����!�z��&���-�����?������g�zi�vJ�$ݰ����M��3�W���b�cd�q�&%M���>"k/;ۃc&i��닕��<L�%�q�ԋ��b}�7�I�%^%ә����*���������B1��:��(�k؍s:��q���%A~��ky񊰞1uf�U	?�S05;�B.��G�B퐂������Px!F��0F<g{�ܓZI�n�!Td�n:;��t��gU�ξ�:=����!C0�A���pã1�y*`��!����~z��}sb��I�{�OB�i��`ȥςT�~�"�v��V�W�@�XlxVHYEB    4ba0    1230��,�!��'�?�,��ǿ�2����Vq��~�|䱍gXg`�+�6HP`����kV����F��9yt��(r���7'D��*x�6���v�D�`�?�D}d�3By�����`��$J(֍���O����d�,�5քĶt\Y "�[�KWyr �}�J¯���5�;�
F�Ơ
�1(r��%��8+��)d\��n�/NXL6�Y�5�	H7�f?�m3x1�V����d��g<`/��A��j��F#�}�� �5��O76���>e�]"�p�7���ٝ�n{�9�2V�U��7����D���[�Q�#�.�_�����\��| {!��<������4�'�.e����ʲ����u'������~MM=�K�҈�X)d=�*��KL��=-B��u��3EI�`s�En���ڀ΃y�7�X�~i��&@� ��[b7,���F�������T�?˟5�k��8ba��I�Sl��|�߅.�ZJbg爰������>�Cj$�]Ū�����,\2h
k$5�۶B���17��������V�˥"W�
��e��A�(qv9�Y���`�������>�5$U})��s�� r�t�#]�/I���IE�qҷO��_<�/���f�Pt���r�.77�q�*�u��@�o1��t�Ļ�4/�,�z����yz>%3';/�(y�~2;V��)����.LV���O��WP�����QH�OgE��;������D�:>t�,��,)Xe]�����2�d��=���`G��^�T� :�v��3D�&�����B_��c��,����u�$Y����bCp�Y7U*|N,ɯ�po�}��?�H/'�t&{MA*	��n0&���7@8��+� z�����܋@N�@����c��o��.��h���ZN�-�`.O��A/����q�e�/��r`�x&��3�>�8�a����xt�*����<Ec�q�	���S�c��H��줨p|s"���I�
ɭM ���k��Nf��'e]X���zM�i w�]J+;�w��N�JW�X���ţ��$�a���4��f�N{��)bgm,E��/��u)� �+��� ��n�u��I�B�D�;6C�$sY�,l��9N[��:�\�qbN�+����Wf�O�_�����q�=hǧ���d˵V�(�}e����/ظ���p���b�ƕ���͉�vQ*�#T�/�5�ˮ�=Y���o<��$����d��\��o�\�8#6�g�8S[䙐�@��������;3����
@I��t�$�Ok�U�n#A�aW�����H��
�
8���s�S�]�%���� �w�:o|�Q�
��L���#̬)��=��x��&7P3�`��M��u�/q�f���J�b־#C_r_�����B����Y�b09}��gn]��D9|�������J�H��UGKlib�k>zh��k�;0U�N�҃�"m�=��`㰬Z���3s�!՜�@ k��u!����Ʃ������U�;�	������GY~��i�Np�Fbe,��+$��FBo�6����;����c>�Y�	�Ǔ"��mD�Y��~a��L�$����bm|_Z[����Qz��r���]��`��"$���`���X��!�7ÕK��Ԓgt��N�� R�Я��-jSj��G2!�j�9K ���2!8
��
��Z�օe<���i��jG�k�tӄ��=悟�OZs�EX�;�zhI&|l�%�`�i�%�?������?�z�+lX��X���D��j� ���*r(Hm�Vm������&82�{�yK��͘�r]�KH����{�6^'�R�;U7��m�>7�)��AL2y)v�s��?޽,d`�y����ou	�
t8y)��dkw��T2��MPl�`x�Ǖ��9@��s��l�?�T-��$�>�M|(��"C$?w�avp6��F�bc���i�5>c�����}^xb����fs-G+�b��]�1�����YI�.Ni:�a�3%(��\P�����p�l���'l��}�Յv�I��vW�>)��h��f�P�(�W��#Ӡ�0!���{����R+ ���%���j?TsE-��[Ղ�f�/BY�ŘO��'�iV����ƫR�Ym�<a	�N�5�r?��1TB����+Uy'":�Z��shO}���i+	#D�����8�D+���������'/(nE��B��8����ė�+�U[m���2���{Z�u��]����f֏&'�8)QA��waY�I��sI����8u������~�-<"u=�kuLW�$MǻIt���Jƹ�]P� �Ԣ�5�r��}f5�V�7����mԒ`欏䷮�ZЗ+QQV��u��KW���/�X�W"Zv���5(-d���
[/�����HQ�[-� �1���	����l�s3k'� ��+Dz���|bCE���EO;O\��;��T��Ma`��Rhb�� ��_��k>'���w�o��o���` eAg�9�6�2�1���gChT�L��NI��v��=(1�NC�V���hg�$%
U4�2��I��Cn�ǘX�����,�Ǣ�-����^H��k�R㇞w�'#a��(�*��L������bi������]��.5�=�=�ꖀ[�G�M�+-�	�u��TE>��SjQ �i�9���	{e�!p:�&��8���l1pͺ�ܵ��h�� �S՜�^PO�B�7���/[al��A)��h�o+i�*�5%�:hę��1V��p��_�ӛ�#bv'��zS�uz��.�m�з���BbY�c�q�?m�gBxWh�
�<b�߅y���_u���Ŀ�K�&�ָs��H��uQ�;֚��j'4�*��e�S�4��\�<A!1��۲|9��쭩���#8�ut��!�ݗ��N.|���Õ:X$�v �|�3ꨄ���H��K�(hS�K��3;bH����Bl�P�{�AJ�Ccg������Ԗͳ�+;���)6�!�����%?�	��?V�fܰك�f�] "ŐEP#��	~��o8Nl	�XtD{�e��S���;���@Һ���{3]}I+��	�M�S��;��O�s?|���[kq�(�k9A0�l�d�4~Fh�Lh��t�*�V=��Rl3�_>0)gǝ�ֳ��6�>�7$�N�n㌩5����;:[/c�Rt�m+�L�a{��'��/�E��z��v�H<���? gn#=k>y˖ӍX���� H2h�W�`=�f��h�c>���O"�H�#�;6H��0"���j�v�-��]b��!���! Mn*���f*"�0⺰g�ɄnD�Gn�0MaN �Ei�f�{�U�4FI���
܃��ݓ��1�_��K�%��}Vf#NN~��l:?Ċ4�O�3���!�G�6���3S^
�!KH���z����@��8\e�.���n�0�ql�tg�VGb����~��3�rq� ��8(S�_)�\c�_�5�v��nn'�^�}2��8��"^�(cέ��RyL�u{qC}� D�)��I�bn3ݤf{O5��Ut[/W�=�(�C�a=F�*��iP7_����j�U�:��t�my}��!+���~������$�� 0"�{mP�%�d<�ُ�("���/O�:����;�(e�Ef�5�r���7�4��bq��K+=Mp�u���D��8w��j����*;�eI�r��X�_j��gx>Hw��1�.2���W�~>u��*=��'�߉Zî�ƌ��b�)v��"r�
�a�m�����k��N�]��+��W��4C5�!���%�5&�	U����] �W�sEΚٽ�wFjx7�#_�	8����%�5x�is}7	�P�*�բ�2�q�2[�t�k9�4C*T@�q,�����2_�u�NT���E�H�?���A;l�DS��V9�/H���H C��#}��9�9
��¾�W��&Q��@@7U�U��4������+�Z�XP�Oԛ��g"�sy.[�܌O.(F����g��E0��N��l���g^�`'�i`#6����l�qa?�kﯯ��o�@k�C�n�J��� T��Z��]�Nt�� ��"峸b
�E�o��/¢+@Y��-�I����3u!s.�r��Tp��m�Lm�s���D$�&B��L�"�d<ґ�[��3�j����՚�%�8�w�KqՍ*}�j�:��\b�RGW��j2���[`V��r½�_8G�J-�Yn���:ȝ����=�z�������|ԣ4�V����}�vR�=�^v�ؖ�N��0���1�Z,�S/�S���Z�o�����2�e�+G�F�,:=-q?m��ȉ����]H��&����"��/�Z��q(_>�ʝ��t���ĥ�v�+�g�\G�f�G6��6I���pw�kw�Rc�h��&X�e1�!�dA�$�ù�h�v�Z��^�}E�����]�/�Ϸ��֪v�p���	8���
z �Qz�`hn?�]����So���Xz`���^�a��|�Fk]-!/km� usf���\
���_�o�z�����'᫐V���[=���hAҖ��