XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��pf�ߢ��kgD�51�Jj�Wp~��N���?!��]�f�L,o0
���1}X|�>t�i���u�5���#��>���Z���Z����7V3_�� xI����Fo88��~�9p����a��
��Ff��b{_�N��w嬣����>��S�,:�jO4Rf:b��3�Ǭϩ�r���r2,�Q+��W��Y�p�Jx{����}�k$��
vm�.?�xw���("�lt�C��-v-�ĩ.x����ӓ��S8��s���
�|xI3?�����NP��#�g_?�oG)S��1��+s�*��k��?�G���X�q6�s}ռ ��y`��N��D�{��uɒ���������X��B�5<ԧɋ�y�-�%xX��]�g�.ă����dߊ�m���D8K���$:�\�ah����!pT����ۃl/`�"D�����엸Ѭn{b�����j�c���v�U�Ч6�|�a:�Eӱ���1ן�n>��n나�T����OU��],$M:�l3#����r':�^�$ԝ�G�8DIX�W�؇O�K}�m]�l )���iGi�@��Ox��=D��� o-\A������������cKl,�/�c�~!z�;Yi^{:Z\J� 4KZ���w�L6���{�fI���w�I^�{�i&��.�xx���t0��@������%��A�:��uv�A<ݿ�W�_��E?�"��`��I�k����5���d����Q�w�����R
�胢�&{	��XlxVHYEB    2bba     bb0H�m�Nr��ž����ܽ��T�/���H�g[y�]:�Y��檏
��)}�E��#�X��2\���S�|PGD��H����w�g^�T?Ҵ��ø\u�:��.�T��i\��:ۼ��
��|�n�!-�.��hv_�a��j6�R�-�@��Ap�W}��J^cc� l�W��e�l������F����n�G!�� ��.lU;;�,�&�X$Y���.aN��ѥ�u��N�tR&�"ۨ�۪!��I[ƣ�8�����~$��;�;4����Êq����,o#`lv��[�&��Z���Ec��;E"��6�#��$��Jir���P��:\yK����)ۆ ��`��� ��\yZ���z� ��WPZ�\a�4 B0PmǷ���w�B
��>���/�߆H��%�}#���]�@���,��OMͪ�=T3�'��D�#Ϙ�;�z�쒱�����`ޑ�����,;kD�5f�|xw�#̮�\WW�c�*R9���w�<k��vO>�s*$%��*+��=m,aF7z`�g��{�RF�T焵m�<+M�BD��u�g�;pe��ܙb��?��n>�8�{V`Z_�b�^�`\t�k�����n��i`����
 }V��HP|�0rP>�ϰK$>v���=�_���R 	(X���	"�S���		M���&�}�"��jUhc��Z�Dc��Fs�*�㫞\@5P��H9������O\���seU��LO�'l#���7H�)[� �E��R���H�&�eF��y�,�s��4�n��'[�<�H��S���7�= Ţ�I�2�R/T�I��U�"���@}H�)��pS�r�f�Ҡ$�{U�_��7$q01�To�X�����I��z�}?��'�P�5��V�H�+Y�8�6M�[X�E��ڡ\�䰠�-�L��%ʛ7c�4���̨��"W8��-�����䛘��H��8j�
�oۍ��͋�i���e�h�zH�������;L�eT�վܩ}`qs*��؀�����u=�9*k<�W�=On�Z
9��խGwT.у�����m(~�Д�\Zh�����z�,��Ǒ���4���s�ľw���c����Z�%�tݐ6O��_�%���{��za�gϣ�32U��� �I�����Č����J�ˑu?�3Ab������#Q������"
9����u�����ޑ�[r�O�
=T��Ju�`��ị�)��`c��u��g��}Ì�|Ɓ�&sE�(��98����>B��׌� q��Ԯ��t#ǽ��ͅA���`�A�g�s�`	�_��^���*��w9k�iX\�E�+_jxYؑ|#ے��&f+_�����OC�����m�S�2'T���vK��W�oP��aH�� }�@yeՆ}�_��E��`;����ǿ� �/5��%�l��bF'*Ö�#[t��&������J-իO���h�uX��T
M���	5ݏ�0�Z���9%�a�Aq:`Ys�Ӵ�_-�T�6b����AuI��������'�sk�0���f�2�c��H��zu�\�Zz���S��NR�z�y<l������}& ��`՞; ��[c�7E~���$\k&�P��y����ƟaUZ�4���%j�4K>u��w@9Q�wL"�2�Ʌ��#Պ��vKD���61�V��o�-Nh�<nМ����,��i��rs��m}\+ݪvuB1ܥ;̬�6X9F�^�L_�`$�#�#ns�^���q��R*�n�����̆ś�HP��$�#���tB����z��ORH���S�'������w�h�|}�3~�(ǘQN9	Y�y?*.b��p���Q�*��[B�c.yG�f���!�zu1�Rs��yX�u�����2&����9p��0��؄���F��ypr�58/��b���c -?|�rF��3���L�ڑ��N�U�.�H_��v�=�5����b?h��3w5�W-��ړ_��Q�A�'��M4so�7��V�1��%��o���(������&���#CH�xh�	~���*����|b�rƐ�yy�'|5!m/h>`M�ҭ���d�i�A3C]��0�~2 �$6�'mX�y���I?�a��K�tE�a��&��N�Ŷ-@1�z��Y�J��Rk�X���+�%��UO��t/��Q	qٚU*ø4tIq��g.��N�b%ؓ:،�7,^��f��ǚR��,� e0�"UbС̐'��b��$|C�yc7'�_0�����b�3��\m�-�\���4�w�&̢>��%�'�TeMi�<����we�1��HOY���h����p�}.�$��e�ª��H�@߈�o�M>C^��:�H�==}B-F����B��ŝ������n�� �I�miz
�)O����eS���V�����w��j�~WnrO�9o������z/�R>c6�^���L	���2�<���:� $�ۨ��S��W7��V]��BHذ�z�_<ݼ��$�|*�1Ζ0>���A�m'������8�G̼�vZ�� F[,ո��s`٠#<��/Ke�HFf司R��Vr`4"}��*&�=��@l�<�����0�jF��"9�2	���@P5�"� ��}�o��3Q����{2�����?{�����HfN"����jRu���e���\)��l����6���.D�Q +B4
����D7Z��Q�oj-(e�D�h�u���9RN���'�~a3����#2P����.;���O�n���s�������/sq�躴������.��R�b�U�?���d������{�g⸾spyYT~5�ts�M�z=�s�Y�>XC|)��1��H�ъw+�aB�>��F��p=�����U�r8�-]��@hJ*H�Mc\�W�������A�4�Z�3��#&D#�ULt������.��2�L[=